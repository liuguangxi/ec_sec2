//==============================================================================
// sect233k1_pt_mul_wrapper.v
//
// Wrapper of module sect233k1_pt_mul.
//------------------------------------------------------------------------------
// Copyright (c) 2022 Guangxi Liu
//
// This source code is licensed under the MIT license found in the
// LICENSE file in the root directory of this source tree.
//==============================================================================


module sect233k1_pt_mul_wrapper (
    // System signals
    input clk,                      // system clock
    input test_i,                   // test input
    output test_o                   // test output
);

// Local signals
wire rst_n;                         // input pin
wire clr;                           // input pin
wire start;                         // input pin
wire [232:0] d;                     // input pin
wire done;                          // output pin
wire [232:0] x;                     // output pin
wire [232:0] y;                     // output pin
wire [235:0] word_o;
wire [466:0] word_i;


// Assignments
assign {rst_n, clr, start, d} = word_o;
assign word_i = {done, x, y};


// Instances
Synthesis_Harness_Input #(
    .WORD_WIDTH     (236)
) u_shi (
    .clock          (clk),
    .clear          (1'b0),
    .bit_in         (test_i),
    .bit_in_valid   (1'b1),
    .word_out       (word_o)
);

Synthesis_Harness_Output #(
    .WORD_WIDTH     (467)
) u_sho (
    .clock          (clk),
    .clear          (1'b0),
    .word_in        (word_i),
    .word_in_valid  (1'b1),
    .bit_out        (test_o)
);

sect233k1_pt_mul u_sect233k1_pt_mul (
    .clk            (clk),
    .rst_n          (rst_n),
    .clr            (clr),
    .start          (start),
    .d              (d),
    .done           (done),
    .x              (x),
    .y              (y)
);


endmodule
